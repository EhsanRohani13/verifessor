module and_testbench;

endmodule
module or_testbench;
initial begin
end
endmodule
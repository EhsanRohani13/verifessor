module and_testbench;
initial begin
end
endmodule